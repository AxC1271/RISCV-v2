`timescale 1ns / 1ps

module hazard_unit (

);

endmodule