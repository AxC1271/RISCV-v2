`timescale 1ns / 1ps

module data_memory (

);

endmodule