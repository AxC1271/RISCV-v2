`timescale 1ns / 1ps

module axi_mmio (
    
);

endmodule