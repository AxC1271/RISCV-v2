`timescale 1ns / 1ps

module instr_cache (

);

endmodule