`timescale 1ns / 1ps

module branch_unit (
    
);

endmodule