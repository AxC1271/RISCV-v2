`timescale 1ns / 1ps

module program_counter (
    input logic clk,
    input logic rst_n,
    input logic[31:0] pc_in,
    output logic[31:0] pc_out
);

endmodule