`timescale 1ns / 1ps;


// derive SVAs for the receiver module
    
module uart_rx_tb();

endmodule